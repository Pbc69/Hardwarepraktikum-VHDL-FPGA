---------------------------------------------------------------------------------------------------
--
-- Titel:    
-- Autor:    
-- Datum:    
-- Laufzeit: 
--
---------------------------------------------------------------------------------------------------

-- Libraries Import:
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
library work;
	use work.all;
	use work.hadescomponents.all;
  
---------------------------------------------------------------------------------------------------

-- Entity:
entity indec_tb is																							   
end indec_tb;																								   
---------------------------------------------------------------------------------------------------


-- Architecture:
architecture TB_ARCHITECTURE of indec_tb is
begin
end TB_ARCHITECTURE;
---------------------------------------------------------------------------------------------------
